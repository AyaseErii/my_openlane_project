VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.720 10.640 30.320 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.080 10.640 45.680 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.440 10.640 61.040 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.800 10.640 76.400 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.160 10.640 91.760 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.520 10.640 107.120 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.400 10.640 38.000 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.760 10.640 53.360 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.120 10.640 68.720 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.480 10.640 84.080 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.200 10.640 114.800 109.040 ;
    END
  END VPWR
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 27.920 120.000 28.520 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 48.320 120.000 48.920 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 50.360 120.000 50.960 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 52.400 120.000 53.000 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 54.440 120.000 55.040 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 56.480 120.000 57.080 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 58.520 120.000 59.120 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 60.560 120.000 61.160 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 62.600 120.000 63.200 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 64.640 120.000 65.240 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 66.680 120.000 67.280 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 29.960 120.000 30.560 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 32.000 120.000 32.600 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 34.040 120.000 34.640 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 36.080 120.000 36.680 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 38.120 120.000 38.720 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 40.160 120.000 40.760 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 42.200 120.000 42.800 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 44.240 120.000 44.840 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 46.280 120.000 46.880 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 68.720 120.000 69.320 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 89.120 120.000 89.720 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 91.160 120.000 91.760 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 93.200 120.000 93.800 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 95.240 120.000 95.840 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 97.280 120.000 97.880 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 99.320 120.000 99.920 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 101.360 120.000 101.960 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 103.400 120.000 104.000 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 105.440 120.000 106.040 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 107.480 120.000 108.080 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 70.760 120.000 71.360 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 72.800 120.000 73.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 74.840 120.000 75.440 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 76.880 120.000 77.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 78.920 120.000 79.520 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 80.960 120.000 81.560 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 83.000 120.000 83.600 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 85.040 120.000 85.640 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 87.080 120.000 87.680 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 116.000 7.730 120.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 116.000 35.330 120.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 116.000 38.090 120.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 116.000 40.850 120.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 116.000 43.610 120.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 116.000 46.370 120.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 116.000 49.130 120.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 116.000 51.890 120.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 116.000 54.650 120.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 116.000 57.410 120.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 116.000 60.170 120.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 116.000 10.490 120.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 116.000 13.250 120.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 116.000 16.010 120.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 116.000 18.770 120.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 116.000 21.530 120.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 116.000 24.290 120.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 116.000 27.050 120.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 116.000 29.810 120.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 116.000 32.570 120.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 116.000 62.930 120.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 116.000 90.530 120.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 116.000 93.290 120.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 116.000 96.050 120.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 116.000 98.810 120.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 116.000 101.570 120.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 116.000 104.330 120.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 116.000 107.090 120.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 116.000 109.850 120.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 116.000 112.610 120.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 116.000 115.370 120.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 116.000 65.690 120.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 116.000 68.450 120.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 116.000 71.210 120.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 116.000 73.970 120.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 116.000 76.730 120.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 116.000 79.490 120.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 116.000 82.250 120.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 116.000 85.010 120.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 116.000 87.770 120.000 ;
    END
  END chany_top_out[9]
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 109.520 120.000 110.120 ;
    END
  END prog_clk_0_E_in
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 19.760 120.000 20.360 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 21.800 120.000 22.400 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 23.840 120.000 24.440 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 25.880 120.000 26.480 ;
    END
  END right_bottom_grid_pin_17_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 9.560 120.000 10.160 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 11.600 120.000 12.200 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 13.640 120.000 14.240 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 15.680 120.000 16.280 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 17.720 120.000 18.320 ;
    END
  END right_bottom_grid_pin_9_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 116.000 4.970 120.000 ;
    END
  END top_left_grid_pin_1_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 4.670 10.640 117.230 109.780 ;
      LAYER met2 ;
        RECT 5.250 115.720 7.170 116.690 ;
        RECT 8.010 115.720 9.930 116.690 ;
        RECT 10.770 115.720 12.690 116.690 ;
        RECT 13.530 115.720 15.450 116.690 ;
        RECT 16.290 115.720 18.210 116.690 ;
        RECT 19.050 115.720 20.970 116.690 ;
        RECT 21.810 115.720 23.730 116.690 ;
        RECT 24.570 115.720 26.490 116.690 ;
        RECT 27.330 115.720 29.250 116.690 ;
        RECT 30.090 115.720 32.010 116.690 ;
        RECT 32.850 115.720 34.770 116.690 ;
        RECT 35.610 115.720 37.530 116.690 ;
        RECT 38.370 115.720 40.290 116.690 ;
        RECT 41.130 115.720 43.050 116.690 ;
        RECT 43.890 115.720 45.810 116.690 ;
        RECT 46.650 115.720 48.570 116.690 ;
        RECT 49.410 115.720 51.330 116.690 ;
        RECT 52.170 115.720 54.090 116.690 ;
        RECT 54.930 115.720 56.850 116.690 ;
        RECT 57.690 115.720 59.610 116.690 ;
        RECT 60.450 115.720 62.370 116.690 ;
        RECT 63.210 115.720 65.130 116.690 ;
        RECT 65.970 115.720 67.890 116.690 ;
        RECT 68.730 115.720 70.650 116.690 ;
        RECT 71.490 115.720 73.410 116.690 ;
        RECT 74.250 115.720 76.170 116.690 ;
        RECT 77.010 115.720 78.930 116.690 ;
        RECT 79.770 115.720 81.690 116.690 ;
        RECT 82.530 115.720 84.450 116.690 ;
        RECT 85.290 115.720 87.210 116.690 ;
        RECT 88.050 115.720 89.970 116.690 ;
        RECT 90.810 115.720 92.730 116.690 ;
        RECT 93.570 115.720 95.490 116.690 ;
        RECT 96.330 115.720 98.250 116.690 ;
        RECT 99.090 115.720 101.010 116.690 ;
        RECT 101.850 115.720 103.770 116.690 ;
        RECT 104.610 115.720 106.530 116.690 ;
        RECT 107.370 115.720 109.290 116.690 ;
        RECT 110.130 115.720 112.050 116.690 ;
        RECT 112.890 115.720 114.810 116.690 ;
        RECT 115.650 115.720 117.200 116.690 ;
        RECT 4.700 9.675 117.200 115.720 ;
      LAYER met3 ;
        RECT 4.000 109.120 115.600 109.985 ;
        RECT 4.000 108.480 116.000 109.120 ;
        RECT 4.000 107.080 115.600 108.480 ;
        RECT 4.000 106.440 116.000 107.080 ;
        RECT 4.000 105.040 115.600 106.440 ;
        RECT 4.000 104.400 116.000 105.040 ;
        RECT 4.000 103.000 115.600 104.400 ;
        RECT 4.000 102.360 116.000 103.000 ;
        RECT 4.000 100.960 115.600 102.360 ;
        RECT 4.000 100.320 116.000 100.960 ;
        RECT 4.000 98.920 115.600 100.320 ;
        RECT 4.000 98.280 116.000 98.920 ;
        RECT 4.000 96.880 115.600 98.280 ;
        RECT 4.000 96.240 116.000 96.880 ;
        RECT 4.000 94.840 115.600 96.240 ;
        RECT 4.000 94.200 116.000 94.840 ;
        RECT 4.000 92.800 115.600 94.200 ;
        RECT 4.000 92.160 116.000 92.800 ;
        RECT 4.000 90.760 115.600 92.160 ;
        RECT 4.000 90.120 116.000 90.760 ;
        RECT 4.400 88.720 115.600 90.120 ;
        RECT 4.000 88.080 116.000 88.720 ;
        RECT 4.000 86.680 115.600 88.080 ;
        RECT 4.000 86.040 116.000 86.680 ;
        RECT 4.000 84.640 115.600 86.040 ;
        RECT 4.000 84.000 116.000 84.640 ;
        RECT 4.000 82.600 115.600 84.000 ;
        RECT 4.000 81.960 116.000 82.600 ;
        RECT 4.000 80.560 115.600 81.960 ;
        RECT 4.000 79.920 116.000 80.560 ;
        RECT 4.000 78.520 115.600 79.920 ;
        RECT 4.000 77.880 116.000 78.520 ;
        RECT 4.000 76.480 115.600 77.880 ;
        RECT 4.000 75.840 116.000 76.480 ;
        RECT 4.000 74.440 115.600 75.840 ;
        RECT 4.000 73.800 116.000 74.440 ;
        RECT 4.000 72.400 115.600 73.800 ;
        RECT 4.000 71.760 116.000 72.400 ;
        RECT 4.000 70.360 115.600 71.760 ;
        RECT 4.000 69.720 116.000 70.360 ;
        RECT 4.000 68.320 115.600 69.720 ;
        RECT 4.000 67.680 116.000 68.320 ;
        RECT 4.000 66.280 115.600 67.680 ;
        RECT 4.000 65.640 116.000 66.280 ;
        RECT 4.000 64.240 115.600 65.640 ;
        RECT 4.000 63.600 116.000 64.240 ;
        RECT 4.000 62.200 115.600 63.600 ;
        RECT 4.000 61.560 116.000 62.200 ;
        RECT 4.000 60.160 115.600 61.560 ;
        RECT 4.000 59.520 116.000 60.160 ;
        RECT 4.000 58.120 115.600 59.520 ;
        RECT 4.000 57.480 116.000 58.120 ;
        RECT 4.000 56.080 115.600 57.480 ;
        RECT 4.000 55.440 116.000 56.080 ;
        RECT 4.000 54.040 115.600 55.440 ;
        RECT 4.000 53.400 116.000 54.040 ;
        RECT 4.000 52.000 115.600 53.400 ;
        RECT 4.000 51.360 116.000 52.000 ;
        RECT 4.000 49.960 115.600 51.360 ;
        RECT 4.000 49.320 116.000 49.960 ;
        RECT 4.000 47.920 115.600 49.320 ;
        RECT 4.000 47.280 116.000 47.920 ;
        RECT 4.000 45.880 115.600 47.280 ;
        RECT 4.000 45.240 116.000 45.880 ;
        RECT 4.000 43.840 115.600 45.240 ;
        RECT 4.000 43.200 116.000 43.840 ;
        RECT 4.000 41.800 115.600 43.200 ;
        RECT 4.000 41.160 116.000 41.800 ;
        RECT 4.000 39.760 115.600 41.160 ;
        RECT 4.000 39.120 116.000 39.760 ;
        RECT 4.000 37.720 115.600 39.120 ;
        RECT 4.000 37.080 116.000 37.720 ;
        RECT 4.000 35.680 115.600 37.080 ;
        RECT 4.000 35.040 116.000 35.680 ;
        RECT 4.000 33.640 115.600 35.040 ;
        RECT 4.000 33.000 116.000 33.640 ;
        RECT 4.000 31.600 115.600 33.000 ;
        RECT 4.000 30.960 116.000 31.600 ;
        RECT 4.000 30.280 115.600 30.960 ;
        RECT 4.400 29.560 115.600 30.280 ;
        RECT 4.400 28.920 116.000 29.560 ;
        RECT 4.400 28.880 115.600 28.920 ;
        RECT 4.000 27.520 115.600 28.880 ;
        RECT 4.000 26.880 116.000 27.520 ;
        RECT 4.000 25.480 115.600 26.880 ;
        RECT 4.000 24.840 116.000 25.480 ;
        RECT 4.000 23.440 115.600 24.840 ;
        RECT 4.000 22.800 116.000 23.440 ;
        RECT 4.000 21.400 115.600 22.800 ;
        RECT 4.000 20.760 116.000 21.400 ;
        RECT 4.000 19.360 115.600 20.760 ;
        RECT 4.000 18.720 116.000 19.360 ;
        RECT 4.000 17.320 115.600 18.720 ;
        RECT 4.000 16.680 116.000 17.320 ;
        RECT 4.000 15.280 115.600 16.680 ;
        RECT 4.000 14.640 116.000 15.280 ;
        RECT 4.000 13.240 115.600 14.640 ;
        RECT 4.000 12.600 116.000 13.240 ;
        RECT 4.000 11.200 115.600 12.600 ;
        RECT 4.000 10.560 116.000 11.200 ;
        RECT 4.000 9.695 115.600 10.560 ;
      LAYER met4 ;
        RECT 103.335 88.575 103.665 104.545 ;
  END
END sb_0__0_
END LIBRARY

