VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__2_
  CLASS BLOCK ;
  FOREIGN sb_0__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 116.000 30.270 120.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END SC_OUT_BOT
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.720 10.640 30.320 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.080 10.640 45.680 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.440 10.640 61.040 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.800 10.640 76.400 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.160 10.640 91.760 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.520 10.640 107.120 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.400 10.640 38.000 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.760 10.640 53.360 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.120 10.640 68.720 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.480 10.640 84.080 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.200 10.640 114.800 109.040 ;
    END
  END VPWR
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END bottom_left_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 116.000 90.070 120.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 25.880 120.000 26.480 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 46.280 120.000 46.880 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 48.320 120.000 48.920 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 50.360 120.000 50.960 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 52.400 120.000 53.000 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 54.440 120.000 55.040 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 56.480 120.000 57.080 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 58.520 120.000 59.120 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 60.560 120.000 61.160 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 62.600 120.000 63.200 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 64.640 120.000 65.240 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 27.920 120.000 28.520 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 29.960 120.000 30.560 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 32.000 120.000 32.600 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 34.040 120.000 34.640 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 36.080 120.000 36.680 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 38.120 120.000 38.720 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 40.160 120.000 40.760 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 42.200 120.000 42.800 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 44.240 120.000 44.840 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 66.680 120.000 67.280 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 87.080 120.000 87.680 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 89.120 120.000 89.720 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 91.160 120.000 91.760 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 93.200 120.000 93.800 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 95.240 120.000 95.840 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 97.280 120.000 97.880 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 99.320 120.000 99.920 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 101.360 120.000 101.960 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 103.400 120.000 104.000 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 105.440 120.000 106.040 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 68.720 120.000 69.320 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 70.760 120.000 71.360 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 72.800 120.000 73.400 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 74.840 120.000 75.440 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 76.880 120.000 77.480 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 78.920 120.000 79.520 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 80.960 120.000 81.560 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 83.000 120.000 83.600 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 85.040 120.000 85.640 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END chany_bottom_out[9]
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 107.480 120.000 108.080 ;
    END
  END prog_clk_0_E_in
  PIN right_bottom_grid_pin_34_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 9.560 120.000 10.160 ;
    END
  END right_bottom_grid_pin_34_
  PIN right_bottom_grid_pin_35_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 11.600 120.000 12.200 ;
    END
  END right_bottom_grid_pin_35_
  PIN right_bottom_grid_pin_36_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 13.640 120.000 14.240 ;
    END
  END right_bottom_grid_pin_36_
  PIN right_bottom_grid_pin_37_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 15.680 120.000 16.280 ;
    END
  END right_bottom_grid_pin_37_
  PIN right_bottom_grid_pin_38_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 17.720 120.000 18.320 ;
    END
  END right_bottom_grid_pin_38_
  PIN right_bottom_grid_pin_39_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 19.760 120.000 20.360 ;
    END
  END right_bottom_grid_pin_39_
  PIN right_bottom_grid_pin_40_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 21.800 120.000 22.400 ;
    END
  END right_bottom_grid_pin_40_
  PIN right_bottom_grid_pin_41_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 23.840 120.000 24.440 ;
    END
  END right_bottom_grid_pin_41_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 109.520 120.000 110.120 ;
    END
  END right_top_grid_pin_1_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 3.290 9.560 116.770 109.040 ;
      LAYER met2 ;
        RECT 3.320 115.720 29.710 116.690 ;
        RECT 30.550 115.720 89.510 116.690 ;
        RECT 90.350 115.720 116.740 116.690 ;
        RECT 3.320 4.280 116.740 115.720 ;
        RECT 3.870 3.670 5.790 4.280 ;
        RECT 6.630 3.670 8.550 4.280 ;
        RECT 9.390 3.670 11.310 4.280 ;
        RECT 12.150 3.670 14.070 4.280 ;
        RECT 14.910 3.670 16.830 4.280 ;
        RECT 17.670 3.670 19.590 4.280 ;
        RECT 20.430 3.670 22.350 4.280 ;
        RECT 23.190 3.670 25.110 4.280 ;
        RECT 25.950 3.670 27.870 4.280 ;
        RECT 28.710 3.670 30.630 4.280 ;
        RECT 31.470 3.670 33.390 4.280 ;
        RECT 34.230 3.670 36.150 4.280 ;
        RECT 36.990 3.670 38.910 4.280 ;
        RECT 39.750 3.670 41.670 4.280 ;
        RECT 42.510 3.670 44.430 4.280 ;
        RECT 45.270 3.670 47.190 4.280 ;
        RECT 48.030 3.670 49.950 4.280 ;
        RECT 50.790 3.670 52.710 4.280 ;
        RECT 53.550 3.670 55.470 4.280 ;
        RECT 56.310 3.670 58.230 4.280 ;
        RECT 59.070 3.670 60.990 4.280 ;
        RECT 61.830 3.670 63.750 4.280 ;
        RECT 64.590 3.670 66.510 4.280 ;
        RECT 67.350 3.670 69.270 4.280 ;
        RECT 70.110 3.670 72.030 4.280 ;
        RECT 72.870 3.670 74.790 4.280 ;
        RECT 75.630 3.670 77.550 4.280 ;
        RECT 78.390 3.670 80.310 4.280 ;
        RECT 81.150 3.670 83.070 4.280 ;
        RECT 83.910 3.670 85.830 4.280 ;
        RECT 86.670 3.670 88.590 4.280 ;
        RECT 89.430 3.670 91.350 4.280 ;
        RECT 92.190 3.670 94.110 4.280 ;
        RECT 94.950 3.670 96.870 4.280 ;
        RECT 97.710 3.670 99.630 4.280 ;
        RECT 100.470 3.670 102.390 4.280 ;
        RECT 103.230 3.670 105.150 4.280 ;
        RECT 105.990 3.670 107.910 4.280 ;
        RECT 108.750 3.670 110.670 4.280 ;
        RECT 111.510 3.670 113.430 4.280 ;
        RECT 114.270 3.670 116.190 4.280 ;
      LAYER met3 ;
        RECT 4.000 109.120 115.600 109.985 ;
        RECT 4.000 108.480 116.000 109.120 ;
        RECT 4.000 107.080 115.600 108.480 ;
        RECT 4.000 106.440 116.000 107.080 ;
        RECT 4.000 105.040 115.600 106.440 ;
        RECT 4.000 104.400 116.000 105.040 ;
        RECT 4.000 103.000 115.600 104.400 ;
        RECT 4.000 102.360 116.000 103.000 ;
        RECT 4.000 100.960 115.600 102.360 ;
        RECT 4.000 100.320 116.000 100.960 ;
        RECT 4.000 98.920 115.600 100.320 ;
        RECT 4.000 98.280 116.000 98.920 ;
        RECT 4.000 96.880 115.600 98.280 ;
        RECT 4.000 96.240 116.000 96.880 ;
        RECT 4.000 94.840 115.600 96.240 ;
        RECT 4.000 94.200 116.000 94.840 ;
        RECT 4.000 92.800 115.600 94.200 ;
        RECT 4.000 92.160 116.000 92.800 ;
        RECT 4.000 90.760 115.600 92.160 ;
        RECT 4.000 90.120 116.000 90.760 ;
        RECT 4.000 88.720 115.600 90.120 ;
        RECT 4.000 88.080 116.000 88.720 ;
        RECT 4.000 86.680 115.600 88.080 ;
        RECT 4.000 86.040 116.000 86.680 ;
        RECT 4.000 84.640 115.600 86.040 ;
        RECT 4.000 84.000 116.000 84.640 ;
        RECT 4.000 82.600 115.600 84.000 ;
        RECT 4.000 81.960 116.000 82.600 ;
        RECT 4.000 80.560 115.600 81.960 ;
        RECT 4.000 79.920 116.000 80.560 ;
        RECT 4.000 78.520 115.600 79.920 ;
        RECT 4.000 77.880 116.000 78.520 ;
        RECT 4.000 76.480 115.600 77.880 ;
        RECT 4.000 75.840 116.000 76.480 ;
        RECT 4.000 74.440 115.600 75.840 ;
        RECT 4.000 73.800 116.000 74.440 ;
        RECT 4.000 72.400 115.600 73.800 ;
        RECT 4.000 71.760 116.000 72.400 ;
        RECT 4.000 70.360 115.600 71.760 ;
        RECT 4.000 69.720 116.000 70.360 ;
        RECT 4.000 68.320 115.600 69.720 ;
        RECT 4.000 67.680 116.000 68.320 ;
        RECT 4.000 66.280 115.600 67.680 ;
        RECT 4.000 65.640 116.000 66.280 ;
        RECT 4.000 64.240 115.600 65.640 ;
        RECT 4.000 63.600 116.000 64.240 ;
        RECT 4.000 62.200 115.600 63.600 ;
        RECT 4.000 61.560 116.000 62.200 ;
        RECT 4.000 60.200 115.600 61.560 ;
        RECT 4.400 60.160 115.600 60.200 ;
        RECT 4.400 59.520 116.000 60.160 ;
        RECT 4.400 58.800 115.600 59.520 ;
        RECT 4.000 58.120 115.600 58.800 ;
        RECT 4.000 57.480 116.000 58.120 ;
        RECT 4.000 56.080 115.600 57.480 ;
        RECT 4.000 55.440 116.000 56.080 ;
        RECT 4.000 54.040 115.600 55.440 ;
        RECT 4.000 53.400 116.000 54.040 ;
        RECT 4.000 52.000 115.600 53.400 ;
        RECT 4.000 51.360 116.000 52.000 ;
        RECT 4.000 49.960 115.600 51.360 ;
        RECT 4.000 49.320 116.000 49.960 ;
        RECT 4.000 47.920 115.600 49.320 ;
        RECT 4.000 47.280 116.000 47.920 ;
        RECT 4.000 45.880 115.600 47.280 ;
        RECT 4.000 45.240 116.000 45.880 ;
        RECT 4.000 43.840 115.600 45.240 ;
        RECT 4.000 43.200 116.000 43.840 ;
        RECT 4.000 41.800 115.600 43.200 ;
        RECT 4.000 41.160 116.000 41.800 ;
        RECT 4.000 39.760 115.600 41.160 ;
        RECT 4.000 39.120 116.000 39.760 ;
        RECT 4.000 37.720 115.600 39.120 ;
        RECT 4.000 37.080 116.000 37.720 ;
        RECT 4.000 35.680 115.600 37.080 ;
        RECT 4.000 35.040 116.000 35.680 ;
        RECT 4.000 33.640 115.600 35.040 ;
        RECT 4.000 33.000 116.000 33.640 ;
        RECT 4.000 31.600 115.600 33.000 ;
        RECT 4.000 30.960 116.000 31.600 ;
        RECT 4.000 29.560 115.600 30.960 ;
        RECT 4.000 28.920 116.000 29.560 ;
        RECT 4.000 27.520 115.600 28.920 ;
        RECT 4.000 26.880 116.000 27.520 ;
        RECT 4.000 25.480 115.600 26.880 ;
        RECT 4.000 24.840 116.000 25.480 ;
        RECT 4.000 23.440 115.600 24.840 ;
        RECT 4.000 22.800 116.000 23.440 ;
        RECT 4.000 21.400 115.600 22.800 ;
        RECT 4.000 20.760 116.000 21.400 ;
        RECT 4.000 19.360 115.600 20.760 ;
        RECT 4.000 18.720 116.000 19.360 ;
        RECT 4.000 17.320 115.600 18.720 ;
        RECT 4.000 16.680 116.000 17.320 ;
        RECT 4.000 15.280 115.600 16.680 ;
        RECT 4.000 14.640 116.000 15.280 ;
        RECT 4.000 13.240 115.600 14.640 ;
        RECT 4.000 12.600 116.000 13.240 ;
        RECT 4.000 11.200 115.600 12.600 ;
        RECT 4.000 10.560 116.000 11.200 ;
        RECT 4.000 9.695 115.600 10.560 ;
      LAYER met4 ;
        RECT 100.575 17.175 104.585 62.385 ;
  END
END sb_0__2_
END LIBRARY

