VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__1_
  CLASS BLOCK ;
  FOREIGN cbx_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 110.000 ;
  PIN REGIN_FEEDTHROUGH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END REGIN_FEEDTHROUGH
  PIN REGOUT_FEEDTHROUGH
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END REGOUT_FEEDTHROUGH
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 106.000 11.870 110.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 106.000 33.490 110.000 ;
    END
  END SC_OUT_TOP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.720 10.640 30.320 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.080 10.640 45.680 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.440 10.640 61.040 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.800 10.640 76.400 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.160 10.640 91.760 98.160 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.400 10.640 38.000 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.760 10.640 53.360 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.120 10.640 68.720 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.480 10.640 84.080 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 98.160 ;
    END
  END VPWR
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_11_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END bottom_grid_pin_11_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_13_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END bottom_grid_pin_13_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_15_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END bottom_grid_pin_15_
  PIN bottom_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END bottom_grid_pin_1_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END bottom_grid_pin_3_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END bottom_grid_pin_5_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END bottom_grid_pin_7_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END bottom_grid_pin_8_
  PIN bottom_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END bottom_grid_pin_9_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 9.560 110.000 10.160 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 29.960 110.000 30.560 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 32.000 110.000 32.600 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 34.040 110.000 34.640 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 36.080 110.000 36.680 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 38.120 110.000 38.720 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 40.160 110.000 40.760 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 42.200 110.000 42.800 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 44.240 110.000 44.840 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 46.280 110.000 46.880 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 48.320 110.000 48.920 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 11.600 110.000 12.200 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 13.640 110.000 14.240 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 15.680 110.000 16.280 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 17.720 110.000 18.320 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 19.760 110.000 20.360 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 21.800 110.000 22.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 23.840 110.000 24.440 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 25.880 110.000 26.480 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 27.920 110.000 28.520 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 50.360 110.000 50.960 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 70.760 110.000 71.360 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 72.800 110.000 73.400 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 74.840 110.000 75.440 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 76.880 110.000 77.480 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 78.920 110.000 79.520 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 80.960 110.000 81.560 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 83.000 110.000 83.600 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 85.040 110.000 85.640 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 87.080 110.000 87.680 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 89.120 110.000 89.720 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 52.400 110.000 53.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 54.440 110.000 55.040 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 56.480 110.000 57.080 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 58.520 110.000 59.120 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 60.560 110.000 61.160 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 62.600 110.000 63.200 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 64.640 110.000 65.240 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 66.680 110.000 67.280 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 68.720 110.000 69.320 ;
    END
  END chanx_right_out[9]
  PIN clk_1_N_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 106.000 55.110 110.000 ;
    END
  END clk_1_N_out
  PIN clk_1_S_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END clk_1_S_out
  PIN clk_1_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END clk_1_W_in
  PIN clk_2_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 91.160 110.000 91.760 ;
    END
  END clk_2_E_out
  PIN clk_2_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END clk_2_W_in
  PIN clk_2_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END clk_2_W_out
  PIN clk_3_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 93.200 110.000 93.800 ;
    END
  END clk_3_E_out
  PIN clk_3_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END clk_3_W_in
  PIN clk_3_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END clk_3_W_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 106.000 76.730 110.000 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 106.000 98.350 110.000 ;
    END
  END prog_clk_0_W_out
  PIN prog_clk_1_N_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 95.240 110.000 95.840 ;
    END
  END prog_clk_1_N_out
  PIN prog_clk_1_S_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END prog_clk_1_S_out
  PIN prog_clk_1_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END prog_clk_1_W_in
  PIN prog_clk_2_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 97.280 110.000 97.880 ;
    END
  END prog_clk_2_E_out
  PIN prog_clk_2_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END prog_clk_2_W_in
  PIN prog_clk_2_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END prog_clk_2_W_out
  PIN prog_clk_3_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.000 99.320 110.000 99.920 ;
    END
  END prog_clk_3_E_out
  PIN prog_clk_3_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END prog_clk_3_W_in
  PIN prog_clk_3_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END prog_clk_3_W_out
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 104.420 98.005 ;
      LAYER met1 ;
        RECT 4.210 6.500 105.730 99.580 ;
      LAYER met2 ;
        RECT 4.240 105.720 11.310 107.285 ;
        RECT 12.150 105.720 32.930 107.285 ;
        RECT 33.770 105.720 54.550 107.285 ;
        RECT 55.390 105.720 76.170 107.285 ;
        RECT 77.010 105.720 97.790 107.285 ;
        RECT 98.630 105.720 105.700 107.285 ;
        RECT 4.240 4.280 105.700 105.720 ;
        RECT 4.240 2.875 6.250 4.280 ;
        RECT 7.090 2.875 10.850 4.280 ;
        RECT 11.690 2.875 15.450 4.280 ;
        RECT 16.290 2.875 20.050 4.280 ;
        RECT 20.890 2.875 24.650 4.280 ;
        RECT 25.490 2.875 29.250 4.280 ;
        RECT 30.090 2.875 33.850 4.280 ;
        RECT 34.690 2.875 38.450 4.280 ;
        RECT 39.290 2.875 43.050 4.280 ;
        RECT 43.890 2.875 47.650 4.280 ;
        RECT 48.490 2.875 52.250 4.280 ;
        RECT 53.090 2.875 56.850 4.280 ;
        RECT 57.690 2.875 61.450 4.280 ;
        RECT 62.290 2.875 66.050 4.280 ;
        RECT 66.890 2.875 70.650 4.280 ;
        RECT 71.490 2.875 75.250 4.280 ;
        RECT 76.090 2.875 79.850 4.280 ;
        RECT 80.690 2.875 84.450 4.280 ;
        RECT 85.290 2.875 89.050 4.280 ;
        RECT 89.890 2.875 93.650 4.280 ;
        RECT 94.490 2.875 98.250 4.280 ;
        RECT 99.090 2.875 102.850 4.280 ;
        RECT 103.690 2.875 105.700 4.280 ;
      LAYER met3 ;
        RECT 4.400 106.400 106.000 107.265 ;
        RECT 4.000 105.760 106.000 106.400 ;
        RECT 4.400 104.360 106.000 105.760 ;
        RECT 4.000 103.720 106.000 104.360 ;
        RECT 4.400 102.320 106.000 103.720 ;
        RECT 4.000 101.680 106.000 102.320 ;
        RECT 4.400 100.320 106.000 101.680 ;
        RECT 4.400 100.280 105.600 100.320 ;
        RECT 4.000 99.640 105.600 100.280 ;
        RECT 4.400 98.920 105.600 99.640 ;
        RECT 4.400 98.280 106.000 98.920 ;
        RECT 4.400 98.240 105.600 98.280 ;
        RECT 4.000 97.600 105.600 98.240 ;
        RECT 4.400 96.880 105.600 97.600 ;
        RECT 4.400 96.240 106.000 96.880 ;
        RECT 4.400 96.200 105.600 96.240 ;
        RECT 4.000 95.560 105.600 96.200 ;
        RECT 4.400 94.840 105.600 95.560 ;
        RECT 4.400 94.200 106.000 94.840 ;
        RECT 4.400 94.160 105.600 94.200 ;
        RECT 4.000 93.520 105.600 94.160 ;
        RECT 4.400 92.800 105.600 93.520 ;
        RECT 4.400 92.160 106.000 92.800 ;
        RECT 4.400 92.120 105.600 92.160 ;
        RECT 4.000 91.480 105.600 92.120 ;
        RECT 4.400 90.760 105.600 91.480 ;
        RECT 4.400 90.120 106.000 90.760 ;
        RECT 4.400 90.080 105.600 90.120 ;
        RECT 4.000 89.440 105.600 90.080 ;
        RECT 4.400 88.720 105.600 89.440 ;
        RECT 4.400 88.080 106.000 88.720 ;
        RECT 4.400 88.040 105.600 88.080 ;
        RECT 4.000 87.400 105.600 88.040 ;
        RECT 4.400 86.680 105.600 87.400 ;
        RECT 4.400 86.040 106.000 86.680 ;
        RECT 4.400 86.000 105.600 86.040 ;
        RECT 4.000 85.360 105.600 86.000 ;
        RECT 4.400 84.640 105.600 85.360 ;
        RECT 4.400 84.000 106.000 84.640 ;
        RECT 4.400 83.960 105.600 84.000 ;
        RECT 4.000 83.320 105.600 83.960 ;
        RECT 4.400 82.600 105.600 83.320 ;
        RECT 4.400 81.960 106.000 82.600 ;
        RECT 4.400 81.920 105.600 81.960 ;
        RECT 4.000 81.280 105.600 81.920 ;
        RECT 4.400 80.560 105.600 81.280 ;
        RECT 4.400 79.920 106.000 80.560 ;
        RECT 4.400 79.880 105.600 79.920 ;
        RECT 4.000 79.240 105.600 79.880 ;
        RECT 4.400 78.520 105.600 79.240 ;
        RECT 4.400 77.880 106.000 78.520 ;
        RECT 4.400 77.840 105.600 77.880 ;
        RECT 4.000 77.200 105.600 77.840 ;
        RECT 4.400 76.480 105.600 77.200 ;
        RECT 4.400 75.840 106.000 76.480 ;
        RECT 4.400 75.800 105.600 75.840 ;
        RECT 4.000 75.160 105.600 75.800 ;
        RECT 4.400 74.440 105.600 75.160 ;
        RECT 4.400 73.800 106.000 74.440 ;
        RECT 4.400 73.760 105.600 73.800 ;
        RECT 4.000 73.120 105.600 73.760 ;
        RECT 4.400 72.400 105.600 73.120 ;
        RECT 4.400 71.760 106.000 72.400 ;
        RECT 4.400 71.720 105.600 71.760 ;
        RECT 4.000 71.080 105.600 71.720 ;
        RECT 4.400 70.360 105.600 71.080 ;
        RECT 4.400 69.720 106.000 70.360 ;
        RECT 4.400 69.680 105.600 69.720 ;
        RECT 4.000 69.040 105.600 69.680 ;
        RECT 4.400 68.320 105.600 69.040 ;
        RECT 4.400 67.680 106.000 68.320 ;
        RECT 4.400 67.640 105.600 67.680 ;
        RECT 4.000 67.000 105.600 67.640 ;
        RECT 4.400 66.280 105.600 67.000 ;
        RECT 4.400 65.640 106.000 66.280 ;
        RECT 4.400 65.600 105.600 65.640 ;
        RECT 4.000 64.960 105.600 65.600 ;
        RECT 4.400 64.240 105.600 64.960 ;
        RECT 4.400 63.600 106.000 64.240 ;
        RECT 4.400 63.560 105.600 63.600 ;
        RECT 4.000 62.920 105.600 63.560 ;
        RECT 4.400 62.200 105.600 62.920 ;
        RECT 4.400 61.560 106.000 62.200 ;
        RECT 4.400 61.520 105.600 61.560 ;
        RECT 4.000 60.880 105.600 61.520 ;
        RECT 4.400 60.160 105.600 60.880 ;
        RECT 4.400 59.520 106.000 60.160 ;
        RECT 4.400 59.480 105.600 59.520 ;
        RECT 4.000 58.840 105.600 59.480 ;
        RECT 4.400 58.120 105.600 58.840 ;
        RECT 4.400 57.480 106.000 58.120 ;
        RECT 4.400 57.440 105.600 57.480 ;
        RECT 4.000 56.800 105.600 57.440 ;
        RECT 4.400 56.080 105.600 56.800 ;
        RECT 4.400 55.440 106.000 56.080 ;
        RECT 4.400 55.400 105.600 55.440 ;
        RECT 4.000 54.760 105.600 55.400 ;
        RECT 4.400 54.040 105.600 54.760 ;
        RECT 4.400 53.400 106.000 54.040 ;
        RECT 4.400 53.360 105.600 53.400 ;
        RECT 4.000 52.720 105.600 53.360 ;
        RECT 4.400 52.000 105.600 52.720 ;
        RECT 4.400 51.360 106.000 52.000 ;
        RECT 4.400 51.320 105.600 51.360 ;
        RECT 4.000 50.680 105.600 51.320 ;
        RECT 4.400 49.960 105.600 50.680 ;
        RECT 4.400 49.320 106.000 49.960 ;
        RECT 4.400 49.280 105.600 49.320 ;
        RECT 4.000 48.640 105.600 49.280 ;
        RECT 4.400 47.920 105.600 48.640 ;
        RECT 4.400 47.280 106.000 47.920 ;
        RECT 4.400 47.240 105.600 47.280 ;
        RECT 4.000 46.600 105.600 47.240 ;
        RECT 4.400 45.880 105.600 46.600 ;
        RECT 4.400 45.240 106.000 45.880 ;
        RECT 4.400 45.200 105.600 45.240 ;
        RECT 4.000 44.560 105.600 45.200 ;
        RECT 4.400 43.840 105.600 44.560 ;
        RECT 4.400 43.200 106.000 43.840 ;
        RECT 4.400 43.160 105.600 43.200 ;
        RECT 4.000 42.520 105.600 43.160 ;
        RECT 4.400 41.800 105.600 42.520 ;
        RECT 4.400 41.160 106.000 41.800 ;
        RECT 4.400 41.120 105.600 41.160 ;
        RECT 4.000 40.480 105.600 41.120 ;
        RECT 4.400 39.760 105.600 40.480 ;
        RECT 4.400 39.120 106.000 39.760 ;
        RECT 4.400 39.080 105.600 39.120 ;
        RECT 4.000 38.440 105.600 39.080 ;
        RECT 4.400 37.720 105.600 38.440 ;
        RECT 4.400 37.080 106.000 37.720 ;
        RECT 4.400 37.040 105.600 37.080 ;
        RECT 4.000 36.400 105.600 37.040 ;
        RECT 4.400 35.680 105.600 36.400 ;
        RECT 4.400 35.040 106.000 35.680 ;
        RECT 4.400 35.000 105.600 35.040 ;
        RECT 4.000 34.360 105.600 35.000 ;
        RECT 4.400 33.640 105.600 34.360 ;
        RECT 4.400 33.000 106.000 33.640 ;
        RECT 4.400 32.960 105.600 33.000 ;
        RECT 4.000 32.320 105.600 32.960 ;
        RECT 4.400 31.600 105.600 32.320 ;
        RECT 4.400 30.960 106.000 31.600 ;
        RECT 4.400 30.920 105.600 30.960 ;
        RECT 4.000 30.280 105.600 30.920 ;
        RECT 4.400 29.560 105.600 30.280 ;
        RECT 4.400 28.920 106.000 29.560 ;
        RECT 4.400 28.880 105.600 28.920 ;
        RECT 4.000 28.240 105.600 28.880 ;
        RECT 4.400 27.520 105.600 28.240 ;
        RECT 4.400 26.880 106.000 27.520 ;
        RECT 4.400 26.840 105.600 26.880 ;
        RECT 4.000 26.200 105.600 26.840 ;
        RECT 4.400 25.480 105.600 26.200 ;
        RECT 4.400 24.840 106.000 25.480 ;
        RECT 4.400 24.800 105.600 24.840 ;
        RECT 4.000 24.160 105.600 24.800 ;
        RECT 4.400 23.440 105.600 24.160 ;
        RECT 4.400 22.800 106.000 23.440 ;
        RECT 4.400 22.760 105.600 22.800 ;
        RECT 4.000 22.120 105.600 22.760 ;
        RECT 4.400 21.400 105.600 22.120 ;
        RECT 4.400 20.760 106.000 21.400 ;
        RECT 4.400 20.720 105.600 20.760 ;
        RECT 4.000 20.080 105.600 20.720 ;
        RECT 4.400 19.360 105.600 20.080 ;
        RECT 4.400 18.720 106.000 19.360 ;
        RECT 4.400 18.680 105.600 18.720 ;
        RECT 4.000 18.040 105.600 18.680 ;
        RECT 4.400 17.320 105.600 18.040 ;
        RECT 4.400 16.680 106.000 17.320 ;
        RECT 4.400 16.640 105.600 16.680 ;
        RECT 4.000 16.000 105.600 16.640 ;
        RECT 4.400 15.280 105.600 16.000 ;
        RECT 4.400 14.640 106.000 15.280 ;
        RECT 4.400 14.600 105.600 14.640 ;
        RECT 4.000 13.960 105.600 14.600 ;
        RECT 4.400 13.240 105.600 13.960 ;
        RECT 4.400 12.600 106.000 13.240 ;
        RECT 4.400 12.560 105.600 12.600 ;
        RECT 4.000 11.920 105.600 12.560 ;
        RECT 4.400 11.200 105.600 11.920 ;
        RECT 4.400 10.560 106.000 11.200 ;
        RECT 4.400 10.520 105.600 10.560 ;
        RECT 4.000 9.880 105.600 10.520 ;
        RECT 4.400 9.160 105.600 9.880 ;
        RECT 4.400 8.480 106.000 9.160 ;
        RECT 4.000 7.840 106.000 8.480 ;
        RECT 4.400 6.440 106.000 7.840 ;
        RECT 4.000 5.800 106.000 6.440 ;
        RECT 4.400 4.400 106.000 5.800 ;
        RECT 4.000 3.760 106.000 4.400 ;
        RECT 4.400 2.895 106.000 3.760 ;
      LAYER met4 ;
        RECT 16.855 11.735 20.640 76.665 ;
        RECT 23.040 11.735 28.320 76.665 ;
        RECT 30.720 11.735 36.000 76.665 ;
        RECT 38.400 11.735 43.680 76.665 ;
        RECT 46.080 11.735 51.360 76.665 ;
        RECT 53.760 11.735 59.040 76.665 ;
        RECT 61.440 11.735 66.720 76.665 ;
        RECT 69.120 11.735 74.400 76.665 ;
        RECT 76.800 11.735 82.080 76.665 ;
        RECT 84.480 11.735 89.760 76.665 ;
        RECT 92.160 11.735 97.225 76.665 ;
  END
END cbx_1__1_
END LIBRARY

