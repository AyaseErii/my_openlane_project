VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 136.000 97.430 140.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 136.000 101.110 140.000 ;
    END
  END SC_OUT_TOP
  PIN Test_en_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 42.200 140.000 42.800 ;
    END
  END Test_en_E_in
  PIN Test_en_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 38.800 140.000 39.400 ;
    END
  END Test_en_E_out
  PIN Test_en_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END Test_en_W_in
  PIN Test_en_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END Test_en_W_out
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.720 10.640 30.320 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.080 10.640 45.680 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.440 10.640 61.040 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.800 10.640 76.400 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.160 10.640 91.760 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.520 10.640 107.120 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.880 10.640 122.480 128.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.400 10.640 38.000 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.760 10.640 53.360 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.120 10.640 68.720 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.480 10.640 84.080 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.200 10.640 114.800 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.560 10.640 130.160 128.080 ;
    END
  END VPWR
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 35.400 140.000 36.000 ;
    END
  END ccff_tail
  PIN clk_0_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 136.000 104.790 140.000 ;
    END
  END clk_0_N_in
  PIN clk_0_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END clk_0_S_in
  PIN prog_clk_0_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 49.000 140.000 49.600 ;
    END
  END prog_clk_0_E_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 45.600 140.000 46.200 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 136.000 108.470 140.000 ;
    END
  END prog_clk_0_N_out
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END prog_clk_0_S_in
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END prog_clk_0_W_out
  PIN right_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 52.400 140.000 53.000 ;
    END
  END right_width_0_height_0__pin_16_
  PIN right_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 55.800 140.000 56.400 ;
    END
  END right_width_0_height_0__pin_17_
  PIN right_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 59.200 140.000 59.800 ;
    END
  END right_width_0_height_0__pin_18_
  PIN right_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 62.600 140.000 63.200 ;
    END
  END right_width_0_height_0__pin_19_
  PIN right_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 66.000 140.000 66.600 ;
    END
  END right_width_0_height_0__pin_20_
  PIN right_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 69.400 140.000 70.000 ;
    END
  END right_width_0_height_0__pin_21_
  PIN right_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 72.800 140.000 73.400 ;
    END
  END right_width_0_height_0__pin_22_
  PIN right_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 76.200 140.000 76.800 ;
    END
  END right_width_0_height_0__pin_23_
  PIN right_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 79.600 140.000 80.200 ;
    END
  END right_width_0_height_0__pin_24_
  PIN right_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 83.000 140.000 83.600 ;
    END
  END right_width_0_height_0__pin_25_
  PIN right_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 86.400 140.000 87.000 ;
    END
  END right_width_0_height_0__pin_26_
  PIN right_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 89.800 140.000 90.400 ;
    END
  END right_width_0_height_0__pin_27_
  PIN right_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 93.200 140.000 93.800 ;
    END
  END right_width_0_height_0__pin_28_
  PIN right_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 96.600 140.000 97.200 ;
    END
  END right_width_0_height_0__pin_29_
  PIN right_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 100.000 140.000 100.600 ;
    END
  END right_width_0_height_0__pin_30_
  PIN right_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 103.400 140.000 104.000 ;
    END
  END right_width_0_height_0__pin_31_
  PIN right_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 8.200 140.000 8.800 ;
    END
  END right_width_0_height_0__pin_42_lower
  PIN right_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 106.800 140.000 107.400 ;
    END
  END right_width_0_height_0__pin_42_upper
  PIN right_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 11.600 140.000 12.200 ;
    END
  END right_width_0_height_0__pin_43_lower
  PIN right_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 110.200 140.000 110.800 ;
    END
  END right_width_0_height_0__pin_43_upper
  PIN right_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 15.000 140.000 15.600 ;
    END
  END right_width_0_height_0__pin_44_lower
  PIN right_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 113.600 140.000 114.200 ;
    END
  END right_width_0_height_0__pin_44_upper
  PIN right_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 18.400 140.000 19.000 ;
    END
  END right_width_0_height_0__pin_45_lower
  PIN right_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 117.000 140.000 117.600 ;
    END
  END right_width_0_height_0__pin_45_upper
  PIN right_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 21.800 140.000 22.400 ;
    END
  END right_width_0_height_0__pin_46_lower
  PIN right_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 120.400 140.000 121.000 ;
    END
  END right_width_0_height_0__pin_46_upper
  PIN right_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 25.200 140.000 25.800 ;
    END
  END right_width_0_height_0__pin_47_lower
  PIN right_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 123.800 140.000 124.400 ;
    END
  END right_width_0_height_0__pin_47_upper
  PIN right_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 28.600 140.000 29.200 ;
    END
  END right_width_0_height_0__pin_48_lower
  PIN right_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 127.200 140.000 127.800 ;
    END
  END right_width_0_height_0__pin_48_upper
  PIN right_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 32.000 140.000 32.600 ;
    END
  END right_width_0_height_0__pin_49_lower
  PIN right_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.000 130.600 140.000 131.200 ;
    END
  END right_width_0_height_0__pin_49_upper
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 136.000 31.190 140.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 136.000 67.990 140.000 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 136.000 71.670 140.000 ;
    END
  END top_width_0_height_0__pin_11_
  PIN top_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 136.000 75.350 140.000 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 136.000 79.030 140.000 ;
    END
  END top_width_0_height_0__pin_13_
  PIN top_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 136.000 82.710 140.000 ;
    END
  END top_width_0_height_0__pin_14_
  PIN top_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 136.000 86.390 140.000 ;
    END
  END top_width_0_height_0__pin_15_
  PIN top_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 136.000 34.870 140.000 ;
    END
  END top_width_0_height_0__pin_1_
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 136.000 38.550 140.000 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 136.000 90.070 140.000 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 136.000 93.750 140.000 ;
    END
  END top_width_0_height_0__pin_33_
  PIN top_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 136.000 112.150 140.000 ;
    END
  END top_width_0_height_0__pin_34_lower
  PIN top_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 136.000 1.750 140.000 ;
    END
  END top_width_0_height_0__pin_34_upper
  PIN top_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 136.000 115.830 140.000 ;
    END
  END top_width_0_height_0__pin_35_lower
  PIN top_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 136.000 5.430 140.000 ;
    END
  END top_width_0_height_0__pin_35_upper
  PIN top_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 136.000 119.510 140.000 ;
    END
  END top_width_0_height_0__pin_36_lower
  PIN top_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 136.000 9.110 140.000 ;
    END
  END top_width_0_height_0__pin_36_upper
  PIN top_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 136.000 123.190 140.000 ;
    END
  END top_width_0_height_0__pin_37_lower
  PIN top_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 136.000 12.790 140.000 ;
    END
  END top_width_0_height_0__pin_37_upper
  PIN top_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 136.000 126.870 140.000 ;
    END
  END top_width_0_height_0__pin_38_lower
  PIN top_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 136.000 16.470 140.000 ;
    END
  END top_width_0_height_0__pin_38_upper
  PIN top_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 136.000 130.550 140.000 ;
    END
  END top_width_0_height_0__pin_39_lower
  PIN top_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 136.000 20.150 140.000 ;
    END
  END top_width_0_height_0__pin_39_upper
  PIN top_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 136.000 42.230 140.000 ;
    END
  END top_width_0_height_0__pin_3_
  PIN top_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 136.000 134.230 140.000 ;
    END
  END top_width_0_height_0__pin_40_lower
  PIN top_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 136.000 23.830 140.000 ;
    END
  END top_width_0_height_0__pin_40_upper
  PIN top_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 136.000 137.910 140.000 ;
    END
  END top_width_0_height_0__pin_41_lower
  PIN top_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 136.000 27.510 140.000 ;
    END
  END top_width_0_height_0__pin_41_upper
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 136.000 45.910 140.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 136.000 49.590 140.000 ;
    END
  END top_width_0_height_0__pin_5_
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 136.000 53.270 140.000 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 136.000 56.950 140.000 ;
    END
  END top_width_0_height_0__pin_7_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 136.000 60.630 140.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 136.000 64.310 140.000 ;
    END
  END top_width_0_height_0__pin_9_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 1.450 10.640 137.930 128.820 ;
      LAYER met2 ;
        RECT 2.030 135.720 4.870 136.410 ;
        RECT 5.710 135.720 8.550 136.410 ;
        RECT 9.390 135.720 12.230 136.410 ;
        RECT 13.070 135.720 15.910 136.410 ;
        RECT 16.750 135.720 19.590 136.410 ;
        RECT 20.430 135.720 23.270 136.410 ;
        RECT 24.110 135.720 26.950 136.410 ;
        RECT 27.790 135.720 30.630 136.410 ;
        RECT 31.470 135.720 34.310 136.410 ;
        RECT 35.150 135.720 37.990 136.410 ;
        RECT 38.830 135.720 41.670 136.410 ;
        RECT 42.510 135.720 45.350 136.410 ;
        RECT 46.190 135.720 49.030 136.410 ;
        RECT 49.870 135.720 52.710 136.410 ;
        RECT 53.550 135.720 56.390 136.410 ;
        RECT 57.230 135.720 60.070 136.410 ;
        RECT 60.910 135.720 63.750 136.410 ;
        RECT 64.590 135.720 67.430 136.410 ;
        RECT 68.270 135.720 71.110 136.410 ;
        RECT 71.950 135.720 74.790 136.410 ;
        RECT 75.630 135.720 78.470 136.410 ;
        RECT 79.310 135.720 82.150 136.410 ;
        RECT 82.990 135.720 85.830 136.410 ;
        RECT 86.670 135.720 89.510 136.410 ;
        RECT 90.350 135.720 93.190 136.410 ;
        RECT 94.030 135.720 96.870 136.410 ;
        RECT 97.710 135.720 100.550 136.410 ;
        RECT 101.390 135.720 104.230 136.410 ;
        RECT 105.070 135.720 107.910 136.410 ;
        RECT 108.750 135.720 111.590 136.410 ;
        RECT 112.430 135.720 115.270 136.410 ;
        RECT 116.110 135.720 118.950 136.410 ;
        RECT 119.790 135.720 122.630 136.410 ;
        RECT 123.470 135.720 126.310 136.410 ;
        RECT 127.150 135.720 129.990 136.410 ;
        RECT 130.830 135.720 133.670 136.410 ;
        RECT 134.510 135.720 137.350 136.410 ;
        RECT 1.480 4.280 137.900 135.720 ;
        RECT 1.480 4.000 11.770 4.280 ;
        RECT 12.610 4.000 34.770 4.280 ;
        RECT 35.610 4.000 57.770 4.280 ;
        RECT 58.610 4.000 80.770 4.280 ;
        RECT 81.610 4.000 103.770 4.280 ;
        RECT 104.610 4.000 126.770 4.280 ;
        RECT 127.610 4.000 137.900 4.280 ;
      LAYER met3 ;
        RECT 4.000 130.200 135.600 131.065 ;
        RECT 4.000 128.200 136.000 130.200 ;
        RECT 4.000 126.800 135.600 128.200 ;
        RECT 4.000 124.800 136.000 126.800 ;
        RECT 4.000 123.400 135.600 124.800 ;
        RECT 4.000 122.760 136.000 123.400 ;
        RECT 4.400 121.400 136.000 122.760 ;
        RECT 4.400 121.360 135.600 121.400 ;
        RECT 4.000 120.000 135.600 121.360 ;
        RECT 4.000 118.000 136.000 120.000 ;
        RECT 4.000 116.600 135.600 118.000 ;
        RECT 4.000 114.600 136.000 116.600 ;
        RECT 4.000 113.200 135.600 114.600 ;
        RECT 4.000 111.200 136.000 113.200 ;
        RECT 4.000 109.800 135.600 111.200 ;
        RECT 4.000 107.800 136.000 109.800 ;
        RECT 4.000 106.400 135.600 107.800 ;
        RECT 4.000 104.400 136.000 106.400 ;
        RECT 4.000 103.000 135.600 104.400 ;
        RECT 4.000 101.000 136.000 103.000 ;
        RECT 4.000 99.600 135.600 101.000 ;
        RECT 4.000 97.600 136.000 99.600 ;
        RECT 4.000 96.200 135.600 97.600 ;
        RECT 4.000 94.200 136.000 96.200 ;
        RECT 4.000 92.800 135.600 94.200 ;
        RECT 4.000 90.800 136.000 92.800 ;
        RECT 4.000 89.400 135.600 90.800 ;
        RECT 4.000 88.080 136.000 89.400 ;
        RECT 4.400 87.400 136.000 88.080 ;
        RECT 4.400 86.680 135.600 87.400 ;
        RECT 4.000 86.000 135.600 86.680 ;
        RECT 4.000 84.000 136.000 86.000 ;
        RECT 4.000 82.600 135.600 84.000 ;
        RECT 4.000 80.600 136.000 82.600 ;
        RECT 4.000 79.200 135.600 80.600 ;
        RECT 4.000 77.200 136.000 79.200 ;
        RECT 4.000 75.800 135.600 77.200 ;
        RECT 4.000 73.800 136.000 75.800 ;
        RECT 4.000 72.400 135.600 73.800 ;
        RECT 4.000 70.400 136.000 72.400 ;
        RECT 4.000 69.000 135.600 70.400 ;
        RECT 4.000 67.000 136.000 69.000 ;
        RECT 4.000 65.600 135.600 67.000 ;
        RECT 4.000 63.600 136.000 65.600 ;
        RECT 4.000 62.200 135.600 63.600 ;
        RECT 4.000 60.200 136.000 62.200 ;
        RECT 4.000 58.800 135.600 60.200 ;
        RECT 4.000 56.800 136.000 58.800 ;
        RECT 4.000 55.400 135.600 56.800 ;
        RECT 4.000 53.400 136.000 55.400 ;
        RECT 4.400 52.000 135.600 53.400 ;
        RECT 4.000 50.000 136.000 52.000 ;
        RECT 4.000 48.600 135.600 50.000 ;
        RECT 4.000 46.600 136.000 48.600 ;
        RECT 4.000 45.200 135.600 46.600 ;
        RECT 4.000 43.200 136.000 45.200 ;
        RECT 4.000 41.800 135.600 43.200 ;
        RECT 4.000 39.800 136.000 41.800 ;
        RECT 4.000 38.400 135.600 39.800 ;
        RECT 4.000 36.400 136.000 38.400 ;
        RECT 4.000 35.000 135.600 36.400 ;
        RECT 4.000 33.000 136.000 35.000 ;
        RECT 4.000 31.600 135.600 33.000 ;
        RECT 4.000 29.600 136.000 31.600 ;
        RECT 4.000 28.200 135.600 29.600 ;
        RECT 4.000 26.200 136.000 28.200 ;
        RECT 4.000 24.800 135.600 26.200 ;
        RECT 4.000 22.800 136.000 24.800 ;
        RECT 4.000 21.400 135.600 22.800 ;
        RECT 4.000 19.400 136.000 21.400 ;
        RECT 4.000 18.720 135.600 19.400 ;
        RECT 4.400 18.000 135.600 18.720 ;
        RECT 4.400 17.320 136.000 18.000 ;
        RECT 4.000 16.000 136.000 17.320 ;
        RECT 4.000 14.600 135.600 16.000 ;
        RECT 4.000 12.600 136.000 14.600 ;
        RECT 4.000 11.200 135.600 12.600 ;
        RECT 4.000 9.200 136.000 11.200 ;
        RECT 4.000 8.335 135.600 9.200 ;
      LAYER met4 ;
        RECT 58.255 31.455 59.040 124.945 ;
        RECT 61.440 31.455 66.720 124.945 ;
        RECT 69.120 31.455 74.400 124.945 ;
        RECT 76.800 31.455 82.080 124.945 ;
        RECT 84.480 31.455 89.760 124.945 ;
        RECT 92.160 31.455 97.440 124.945 ;
        RECT 99.840 31.455 105.120 124.945 ;
        RECT 107.520 31.455 112.800 124.945 ;
        RECT 115.200 31.455 120.480 124.945 ;
        RECT 122.880 31.455 127.585 124.945 ;
  END
END grid_clb
END LIBRARY

