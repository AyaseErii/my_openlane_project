VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tie_array
  CLASS BLOCK ;
  FOREIGN tie_array ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 55.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.720 10.640 30.320 54.640 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.400 10.640 38.000 54.640 ;
    END
  END VPWR
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END x[7]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 44.160 54.485 ;
      LAYER met1 ;
        RECT 3.750 10.640 45.930 54.640 ;
      LAYER met2 ;
        RECT 3.780 4.280 45.900 54.585 ;
        RECT 4.330 4.000 9.470 4.280 ;
        RECT 10.310 4.000 15.450 4.280 ;
        RECT 16.290 4.000 21.430 4.280 ;
        RECT 22.270 4.000 27.410 4.280 ;
        RECT 28.250 4.000 33.390 4.280 ;
        RECT 34.230 4.000 39.370 4.280 ;
        RECT 40.210 4.000 45.350 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 37.990 54.565 ;
  END
END tie_array
END LIBRARY

