VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__2_
  CLASS BLOCK ;
  FOREIGN cbx_1__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 210.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 200.000 82.240 ;
    END
  END IO_ISOL_N
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 206.000 71.210 210.000 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 206.000 119.510 210.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END SC_OUT_TOP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 198.800 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 198.800 ;
    END
  END VPWR
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_11_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END bottom_grid_pin_11_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 206.000 61.550 210.000 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_13_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END bottom_grid_pin_13_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_15_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 206.000 177.470 210.000 ;
    END
  END bottom_grid_pin_15_
  PIN bottom_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END bottom_grid_pin_1_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.040 200.000 187.640 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END bottom_grid_pin_3_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 13.640 200.000 14.240 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.040 200.000 170.640 ;
    END
  END bottom_grid_pin_5_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 206.000 96.970 210.000 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 206.000 26.130 210.000 ;
    END
  END bottom_grid_pin_7_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 193.840 200.000 194.440 ;
    END
  END bottom_grid_pin_8_
  PIN bottom_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 206.000 48.670 210.000 ;
    END
  END bottom_grid_pin_9_
  PIN bottom_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END bottom_width_0_height_0__pin_0_
  PIN bottom_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END bottom_width_0_height_0__pin_1_lower
  PIN bottom_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END bottom_width_0_height_0__pin_1_upper
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 206.000 106.630 210.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 206.000 84.090 210.000 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 51.040 200.000 51.640 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 206.000 161.370 210.000 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 57.840 200.000 58.440 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 180.240 200.000 180.840 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 156.440 200.000 157.040 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 142.840 200.000 143.440 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 132.640 200.000 133.240 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 200.640 200.000 201.240 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 206.000 90.530 210.000 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 105.440 200.000 106.040 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 112.240 200.000 112.840 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 206.000 55.110 210.000 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 206.000 113.070 210.000 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 206.000 183.910 210.000 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 44.240 200.000 44.840 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 20.440 200.000 21.040 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 37.440 200.000 38.040 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 206.000 196.790 210.000 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 64.640 200.000 65.240 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 206.000 42.230 210.000 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 6.840 200.000 7.440 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 206.000 135.610 210.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 0.040 200.000 0.640 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.040 200.000 119.640 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 74.840 200.000 75.440 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 88.440 200.000 89.040 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 149.640 200.000 150.240 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 163.240 200.000 163.840 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 206.000 13.250 210.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 206.000 19.690 210.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 206.000 77.650 210.000 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 206.000 142.050 210.000 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 206.000 171.030 210.000 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 206.000 125.950 210.000 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 206.000 190.350 210.000 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 27.240 200.000 27.840 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.840 200.000 126.440 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 206.000 154.930 210.000 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 206.000 148.490 210.000 ;
    END
  END chanx_right_out[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 206.000 6.810 210.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 206.000 35.790 210.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END prog_clk_0_S_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END prog_clk_0_W_out
  PIN top_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 200.000 95.840 ;
    END
  END top_grid_pin_0_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 198.645 ;
      LAYER met1 ;
        RECT 0.070 10.640 196.810 198.800 ;
      LAYER met2 ;
        RECT 0.100 205.720 6.250 207.925 ;
        RECT 7.090 205.720 12.690 207.925 ;
        RECT 13.530 205.720 19.130 207.925 ;
        RECT 19.970 205.720 25.570 207.925 ;
        RECT 26.410 205.720 35.230 207.925 ;
        RECT 36.070 205.720 41.670 207.925 ;
        RECT 42.510 205.720 48.110 207.925 ;
        RECT 48.950 205.720 54.550 207.925 ;
        RECT 55.390 205.720 60.990 207.925 ;
        RECT 61.830 205.720 70.650 207.925 ;
        RECT 71.490 205.720 77.090 207.925 ;
        RECT 77.930 205.720 83.530 207.925 ;
        RECT 84.370 205.720 89.970 207.925 ;
        RECT 90.810 205.720 96.410 207.925 ;
        RECT 97.250 205.720 106.070 207.925 ;
        RECT 106.910 205.720 112.510 207.925 ;
        RECT 113.350 205.720 118.950 207.925 ;
        RECT 119.790 205.720 125.390 207.925 ;
        RECT 126.230 205.720 135.050 207.925 ;
        RECT 135.890 205.720 141.490 207.925 ;
        RECT 142.330 205.720 147.930 207.925 ;
        RECT 148.770 205.720 154.370 207.925 ;
        RECT 155.210 205.720 160.810 207.925 ;
        RECT 161.650 205.720 170.470 207.925 ;
        RECT 171.310 205.720 176.910 207.925 ;
        RECT 177.750 205.720 183.350 207.925 ;
        RECT 184.190 205.720 189.790 207.925 ;
        RECT 190.630 205.720 196.230 207.925 ;
        RECT 0.100 4.280 196.780 205.720 ;
        RECT 0.650 0.155 6.250 4.280 ;
        RECT 7.090 0.155 12.690 4.280 ;
        RECT 13.530 0.155 19.130 4.280 ;
        RECT 19.970 0.155 25.570 4.280 ;
        RECT 26.410 0.155 35.230 4.280 ;
        RECT 36.070 0.155 41.670 4.280 ;
        RECT 42.510 0.155 48.110 4.280 ;
        RECT 48.950 0.155 54.550 4.280 ;
        RECT 55.390 0.155 60.990 4.280 ;
        RECT 61.830 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 83.530 4.280 ;
        RECT 84.370 0.155 89.970 4.280 ;
        RECT 90.810 0.155 99.630 4.280 ;
        RECT 100.470 0.155 106.070 4.280 ;
        RECT 106.910 0.155 112.510 4.280 ;
        RECT 113.350 0.155 118.950 4.280 ;
        RECT 119.790 0.155 125.390 4.280 ;
        RECT 126.230 0.155 135.050 4.280 ;
        RECT 135.890 0.155 141.490 4.280 ;
        RECT 142.330 0.155 147.930 4.280 ;
        RECT 148.770 0.155 154.370 4.280 ;
        RECT 155.210 0.155 160.810 4.280 ;
        RECT 161.650 0.155 170.470 4.280 ;
        RECT 171.310 0.155 176.910 4.280 ;
        RECT 177.750 0.155 183.350 4.280 ;
        RECT 184.190 0.155 189.790 4.280 ;
        RECT 190.630 0.155 196.780 4.280 ;
      LAYER met3 ;
        RECT 4.400 207.040 196.000 207.905 ;
        RECT 4.000 201.640 196.000 207.040 ;
        RECT 4.400 200.240 195.600 201.640 ;
        RECT 4.000 194.840 196.000 200.240 ;
        RECT 4.400 193.440 195.600 194.840 ;
        RECT 4.000 188.040 196.000 193.440 ;
        RECT 4.400 186.640 195.600 188.040 ;
        RECT 4.000 181.240 196.000 186.640 ;
        RECT 4.400 179.840 195.600 181.240 ;
        RECT 4.000 171.040 196.000 179.840 ;
        RECT 4.400 169.640 195.600 171.040 ;
        RECT 4.000 164.240 196.000 169.640 ;
        RECT 4.400 162.840 195.600 164.240 ;
        RECT 4.000 157.440 196.000 162.840 ;
        RECT 4.400 156.040 195.600 157.440 ;
        RECT 4.000 150.640 196.000 156.040 ;
        RECT 4.400 149.240 195.600 150.640 ;
        RECT 4.000 143.840 196.000 149.240 ;
        RECT 4.400 142.440 195.600 143.840 ;
        RECT 4.000 133.640 196.000 142.440 ;
        RECT 4.400 132.240 195.600 133.640 ;
        RECT 4.000 126.840 196.000 132.240 ;
        RECT 4.400 125.440 195.600 126.840 ;
        RECT 4.000 120.040 196.000 125.440 ;
        RECT 4.400 118.640 195.600 120.040 ;
        RECT 4.000 113.240 196.000 118.640 ;
        RECT 4.400 111.840 195.600 113.240 ;
        RECT 4.000 106.440 196.000 111.840 ;
        RECT 4.000 105.040 195.600 106.440 ;
        RECT 4.000 103.040 196.000 105.040 ;
        RECT 4.400 101.640 196.000 103.040 ;
        RECT 4.000 96.240 196.000 101.640 ;
        RECT 4.400 94.840 195.600 96.240 ;
        RECT 4.000 89.440 196.000 94.840 ;
        RECT 4.400 88.040 195.600 89.440 ;
        RECT 4.000 82.640 196.000 88.040 ;
        RECT 4.400 81.240 195.600 82.640 ;
        RECT 4.000 75.840 196.000 81.240 ;
        RECT 4.400 74.440 195.600 75.840 ;
        RECT 4.000 65.640 196.000 74.440 ;
        RECT 4.400 64.240 195.600 65.640 ;
        RECT 4.000 58.840 196.000 64.240 ;
        RECT 4.400 57.440 195.600 58.840 ;
        RECT 4.000 52.040 196.000 57.440 ;
        RECT 4.400 50.640 195.600 52.040 ;
        RECT 4.000 45.240 196.000 50.640 ;
        RECT 4.400 43.840 195.600 45.240 ;
        RECT 4.000 38.440 196.000 43.840 ;
        RECT 4.400 37.040 195.600 38.440 ;
        RECT 4.000 28.240 196.000 37.040 ;
        RECT 4.400 26.840 195.600 28.240 ;
        RECT 4.000 21.440 196.000 26.840 ;
        RECT 4.400 20.040 195.600 21.440 ;
        RECT 4.000 14.640 196.000 20.040 ;
        RECT 4.400 13.240 195.600 14.640 ;
        RECT 4.000 7.840 196.000 13.240 ;
        RECT 4.400 6.440 195.600 7.840 ;
        RECT 4.000 1.040 196.000 6.440 ;
        RECT 4.000 0.175 195.600 1.040 ;
  END
END cbx_1__2_
END LIBRARY

