VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__1_
  CLASS BLOCK ;
  FOREIGN sb_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.720 10.640 30.320 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.080 10.640 45.680 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.440 10.640 61.040 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.800 10.640 76.400 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.160 10.640 91.760 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.520 10.640 107.120 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.400 10.640 38.000 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.760 10.640 53.360 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.120 10.640 68.720 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.480 10.640 84.080 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.200 10.640 114.800 109.040 ;
    END
  END VPWR
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END bottom_left_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 26.560 120.000 27.160 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 46.960 120.000 47.560 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 49.000 120.000 49.600 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 51.040 120.000 51.640 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 53.080 120.000 53.680 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 55.120 120.000 55.720 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 57.160 120.000 57.760 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 59.200 120.000 59.800 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 61.240 120.000 61.840 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 63.280 120.000 63.880 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 65.320 120.000 65.920 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 28.600 120.000 29.200 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 30.640 120.000 31.240 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 32.680 120.000 33.280 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 34.720 120.000 35.320 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 36.760 120.000 37.360 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 38.800 120.000 39.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 40.840 120.000 41.440 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 42.880 120.000 43.480 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 44.920 120.000 45.520 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 67.360 120.000 67.960 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 87.760 120.000 88.360 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 89.800 120.000 90.400 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 91.840 120.000 92.440 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 93.880 120.000 94.480 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 95.920 120.000 96.520 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 97.960 120.000 98.560 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 100.000 120.000 100.600 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 102.040 120.000 102.640 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 104.080 120.000 104.680 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 106.120 120.000 106.720 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 69.400 120.000 70.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 71.440 120.000 72.040 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 73.480 120.000 74.080 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 75.520 120.000 76.120 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 77.560 120.000 78.160 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 79.600 120.000 80.200 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 81.640 120.000 82.240 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 83.680 120.000 84.280 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 85.720 120.000 86.320 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 116.000 7.730 120.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 116.000 35.330 120.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 116.000 38.090 120.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 116.000 40.850 120.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 116.000 43.610 120.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 116.000 46.370 120.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 116.000 49.130 120.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 116.000 51.890 120.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 116.000 54.650 120.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 116.000 57.410 120.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 116.000 60.170 120.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 116.000 10.490 120.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 116.000 13.250 120.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 116.000 16.010 120.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 116.000 18.770 120.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 116.000 21.530 120.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 116.000 24.290 120.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 116.000 27.050 120.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 116.000 29.810 120.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 116.000 32.570 120.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 116.000 62.930 120.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 116.000 90.530 120.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 116.000 93.290 120.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 116.000 96.050 120.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 116.000 98.810 120.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 116.000 101.570 120.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 116.000 104.330 120.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 116.000 107.090 120.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 116.000 109.850 120.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 116.000 112.610 120.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 116.000 115.370 120.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 116.000 65.690 120.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 116.000 68.450 120.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 116.000 71.210 120.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 116.000 73.970 120.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 116.000 76.730 120.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 116.000 79.490 120.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 116.000 82.250 120.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 116.000 85.010 120.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 116.000 87.770 120.000 ;
    END
  END chany_top_out[9]
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 108.160 120.000 108.760 ;
    END
  END prog_clk_0_E_in
  PIN right_bottom_grid_pin_34_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 10.240 120.000 10.840 ;
    END
  END right_bottom_grid_pin_34_
  PIN right_bottom_grid_pin_35_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 12.280 120.000 12.880 ;
    END
  END right_bottom_grid_pin_35_
  PIN right_bottom_grid_pin_36_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 14.320 120.000 14.920 ;
    END
  END right_bottom_grid_pin_36_
  PIN right_bottom_grid_pin_37_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 16.360 120.000 16.960 ;
    END
  END right_bottom_grid_pin_37_
  PIN right_bottom_grid_pin_38_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 18.400 120.000 19.000 ;
    END
  END right_bottom_grid_pin_38_
  PIN right_bottom_grid_pin_39_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 20.440 120.000 21.040 ;
    END
  END right_bottom_grid_pin_39_
  PIN right_bottom_grid_pin_40_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 22.480 120.000 23.080 ;
    END
  END right_bottom_grid_pin_40_
  PIN right_bottom_grid_pin_41_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000 24.520 120.000 25.120 ;
    END
  END right_bottom_grid_pin_41_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 116.000 4.970 120.000 ;
    END
  END top_left_grid_pin_1_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 4.670 10.240 115.390 109.040 ;
      LAYER met2 ;
        RECT 5.250 115.720 7.170 116.690 ;
        RECT 8.010 115.720 9.930 116.690 ;
        RECT 10.770 115.720 12.690 116.690 ;
        RECT 13.530 115.720 15.450 116.690 ;
        RECT 16.290 115.720 18.210 116.690 ;
        RECT 19.050 115.720 20.970 116.690 ;
        RECT 21.810 115.720 23.730 116.690 ;
        RECT 24.570 115.720 26.490 116.690 ;
        RECT 27.330 115.720 29.250 116.690 ;
        RECT 30.090 115.720 32.010 116.690 ;
        RECT 32.850 115.720 34.770 116.690 ;
        RECT 35.610 115.720 37.530 116.690 ;
        RECT 38.370 115.720 40.290 116.690 ;
        RECT 41.130 115.720 43.050 116.690 ;
        RECT 43.890 115.720 45.810 116.690 ;
        RECT 46.650 115.720 48.570 116.690 ;
        RECT 49.410 115.720 51.330 116.690 ;
        RECT 52.170 115.720 54.090 116.690 ;
        RECT 54.930 115.720 56.850 116.690 ;
        RECT 57.690 115.720 59.610 116.690 ;
        RECT 60.450 115.720 62.370 116.690 ;
        RECT 63.210 115.720 65.130 116.690 ;
        RECT 65.970 115.720 67.890 116.690 ;
        RECT 68.730 115.720 70.650 116.690 ;
        RECT 71.490 115.720 73.410 116.690 ;
        RECT 74.250 115.720 76.170 116.690 ;
        RECT 77.010 115.720 78.930 116.690 ;
        RECT 79.770 115.720 81.690 116.690 ;
        RECT 82.530 115.720 84.450 116.690 ;
        RECT 85.290 115.720 87.210 116.690 ;
        RECT 88.050 115.720 89.970 116.690 ;
        RECT 90.810 115.720 92.730 116.690 ;
        RECT 93.570 115.720 95.490 116.690 ;
        RECT 96.330 115.720 98.250 116.690 ;
        RECT 99.090 115.720 101.010 116.690 ;
        RECT 101.850 115.720 103.770 116.690 ;
        RECT 104.610 115.720 106.530 116.690 ;
        RECT 107.370 115.720 109.290 116.690 ;
        RECT 110.130 115.720 112.050 116.690 ;
        RECT 112.890 115.720 114.810 116.690 ;
        RECT 4.700 4.280 115.360 115.720 ;
        RECT 5.250 3.670 7.170 4.280 ;
        RECT 8.010 3.670 9.930 4.280 ;
        RECT 10.770 3.670 12.690 4.280 ;
        RECT 13.530 3.670 15.450 4.280 ;
        RECT 16.290 3.670 18.210 4.280 ;
        RECT 19.050 3.670 20.970 4.280 ;
        RECT 21.810 3.670 23.730 4.280 ;
        RECT 24.570 3.670 26.490 4.280 ;
        RECT 27.330 3.670 29.250 4.280 ;
        RECT 30.090 3.670 32.010 4.280 ;
        RECT 32.850 3.670 34.770 4.280 ;
        RECT 35.610 3.670 37.530 4.280 ;
        RECT 38.370 3.670 40.290 4.280 ;
        RECT 41.130 3.670 43.050 4.280 ;
        RECT 43.890 3.670 45.810 4.280 ;
        RECT 46.650 3.670 48.570 4.280 ;
        RECT 49.410 3.670 51.330 4.280 ;
        RECT 52.170 3.670 54.090 4.280 ;
        RECT 54.930 3.670 56.850 4.280 ;
        RECT 57.690 3.670 59.610 4.280 ;
        RECT 60.450 3.670 62.370 4.280 ;
        RECT 63.210 3.670 65.130 4.280 ;
        RECT 65.970 3.670 67.890 4.280 ;
        RECT 68.730 3.670 70.650 4.280 ;
        RECT 71.490 3.670 73.410 4.280 ;
        RECT 74.250 3.670 76.170 4.280 ;
        RECT 77.010 3.670 78.930 4.280 ;
        RECT 79.770 3.670 81.690 4.280 ;
        RECT 82.530 3.670 84.450 4.280 ;
        RECT 85.290 3.670 87.210 4.280 ;
        RECT 88.050 3.670 89.970 4.280 ;
        RECT 90.810 3.670 92.730 4.280 ;
        RECT 93.570 3.670 95.490 4.280 ;
        RECT 96.330 3.670 98.250 4.280 ;
        RECT 99.090 3.670 101.010 4.280 ;
        RECT 101.850 3.670 103.770 4.280 ;
        RECT 104.610 3.670 106.530 4.280 ;
        RECT 107.370 3.670 109.290 4.280 ;
        RECT 110.130 3.670 112.050 4.280 ;
        RECT 112.890 3.670 114.810 4.280 ;
      LAYER met3 ;
        RECT 4.000 107.760 115.600 108.965 ;
        RECT 4.000 107.120 116.000 107.760 ;
        RECT 4.000 105.720 115.600 107.120 ;
        RECT 4.000 105.080 116.000 105.720 ;
        RECT 4.000 103.680 115.600 105.080 ;
        RECT 4.000 103.040 116.000 103.680 ;
        RECT 4.000 101.640 115.600 103.040 ;
        RECT 4.000 101.000 116.000 101.640 ;
        RECT 4.000 99.600 115.600 101.000 ;
        RECT 4.000 98.960 116.000 99.600 ;
        RECT 4.000 97.560 115.600 98.960 ;
        RECT 4.000 96.920 116.000 97.560 ;
        RECT 4.000 95.520 115.600 96.920 ;
        RECT 4.000 94.880 116.000 95.520 ;
        RECT 4.000 93.480 115.600 94.880 ;
        RECT 4.000 92.840 116.000 93.480 ;
        RECT 4.000 91.440 115.600 92.840 ;
        RECT 4.000 90.800 116.000 91.440 ;
        RECT 4.000 90.120 115.600 90.800 ;
        RECT 4.400 89.400 115.600 90.120 ;
        RECT 4.400 88.760 116.000 89.400 ;
        RECT 4.400 88.720 115.600 88.760 ;
        RECT 4.000 87.360 115.600 88.720 ;
        RECT 4.000 86.720 116.000 87.360 ;
        RECT 4.000 85.320 115.600 86.720 ;
        RECT 4.000 84.680 116.000 85.320 ;
        RECT 4.000 83.280 115.600 84.680 ;
        RECT 4.000 82.640 116.000 83.280 ;
        RECT 4.000 81.240 115.600 82.640 ;
        RECT 4.000 80.600 116.000 81.240 ;
        RECT 4.000 79.200 115.600 80.600 ;
        RECT 4.000 78.560 116.000 79.200 ;
        RECT 4.000 77.160 115.600 78.560 ;
        RECT 4.000 76.520 116.000 77.160 ;
        RECT 4.000 75.120 115.600 76.520 ;
        RECT 4.000 74.480 116.000 75.120 ;
        RECT 4.000 73.080 115.600 74.480 ;
        RECT 4.000 72.440 116.000 73.080 ;
        RECT 4.000 71.040 115.600 72.440 ;
        RECT 4.000 70.400 116.000 71.040 ;
        RECT 4.000 69.000 115.600 70.400 ;
        RECT 4.000 68.360 116.000 69.000 ;
        RECT 4.000 66.960 115.600 68.360 ;
        RECT 4.000 66.320 116.000 66.960 ;
        RECT 4.000 64.920 115.600 66.320 ;
        RECT 4.000 64.280 116.000 64.920 ;
        RECT 4.000 62.880 115.600 64.280 ;
        RECT 4.000 62.240 116.000 62.880 ;
        RECT 4.000 60.840 115.600 62.240 ;
        RECT 4.000 60.200 116.000 60.840 ;
        RECT 4.000 58.800 115.600 60.200 ;
        RECT 4.000 58.160 116.000 58.800 ;
        RECT 4.000 56.760 115.600 58.160 ;
        RECT 4.000 56.120 116.000 56.760 ;
        RECT 4.000 54.720 115.600 56.120 ;
        RECT 4.000 54.080 116.000 54.720 ;
        RECT 4.000 52.680 115.600 54.080 ;
        RECT 4.000 52.040 116.000 52.680 ;
        RECT 4.000 50.640 115.600 52.040 ;
        RECT 4.000 50.000 116.000 50.640 ;
        RECT 4.000 48.600 115.600 50.000 ;
        RECT 4.000 47.960 116.000 48.600 ;
        RECT 4.000 46.560 115.600 47.960 ;
        RECT 4.000 45.920 116.000 46.560 ;
        RECT 4.000 44.520 115.600 45.920 ;
        RECT 4.000 43.880 116.000 44.520 ;
        RECT 4.000 42.480 115.600 43.880 ;
        RECT 4.000 41.840 116.000 42.480 ;
        RECT 4.000 40.440 115.600 41.840 ;
        RECT 4.000 39.800 116.000 40.440 ;
        RECT 4.000 38.400 115.600 39.800 ;
        RECT 4.000 37.760 116.000 38.400 ;
        RECT 4.000 36.360 115.600 37.760 ;
        RECT 4.000 35.720 116.000 36.360 ;
        RECT 4.000 34.320 115.600 35.720 ;
        RECT 4.000 33.680 116.000 34.320 ;
        RECT 4.000 32.280 115.600 33.680 ;
        RECT 4.000 31.640 116.000 32.280 ;
        RECT 4.000 30.280 115.600 31.640 ;
        RECT 4.400 30.240 115.600 30.280 ;
        RECT 4.400 29.600 116.000 30.240 ;
        RECT 4.400 28.880 115.600 29.600 ;
        RECT 4.000 28.200 115.600 28.880 ;
        RECT 4.000 27.560 116.000 28.200 ;
        RECT 4.000 26.160 115.600 27.560 ;
        RECT 4.000 25.520 116.000 26.160 ;
        RECT 4.000 24.120 115.600 25.520 ;
        RECT 4.000 23.480 116.000 24.120 ;
        RECT 4.000 22.080 115.600 23.480 ;
        RECT 4.000 21.440 116.000 22.080 ;
        RECT 4.000 20.040 115.600 21.440 ;
        RECT 4.000 19.400 116.000 20.040 ;
        RECT 4.000 18.000 115.600 19.400 ;
        RECT 4.000 17.360 116.000 18.000 ;
        RECT 4.000 15.960 115.600 17.360 ;
        RECT 4.000 15.320 116.000 15.960 ;
        RECT 4.000 13.920 115.600 15.320 ;
        RECT 4.000 13.280 116.000 13.920 ;
        RECT 4.000 11.880 115.600 13.280 ;
        RECT 4.000 11.240 116.000 11.880 ;
        RECT 4.000 10.390 115.600 11.240 ;
      LAYER met4 ;
        RECT 38.935 11.735 43.680 97.065 ;
        RECT 46.080 11.735 51.360 97.065 ;
        RECT 53.760 11.735 59.040 97.065 ;
        RECT 61.440 11.735 66.720 97.065 ;
        RECT 69.120 11.735 74.400 97.065 ;
        RECT 76.800 11.735 82.080 97.065 ;
        RECT 84.480 11.735 89.760 97.065 ;
        RECT 92.160 11.735 97.440 97.065 ;
        RECT 99.840 11.735 102.745 97.065 ;
  END
END sb_0__1_
END LIBRARY

